module empty;
endmodule